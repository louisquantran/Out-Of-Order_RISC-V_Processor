`timescale 1ns / 1ps

import types_pkg::*;

module fu_mem(
    input clk,
    input reset,
        
    // From ROB
    input logic retired,
    input logic [4:0] rob_head,
    input logic [4:0] curr_rob_tag,
    input logic mispredict,
    input logic [4:0] mispredict_tag,
    
    // From RS and PRF
    input logic issued,
    input rs_data data_in,
    input logic [31:0] ps1_data,
    input logic [31:0] ps2_data,
    
    // Output data
    output mem_data data_out
);
    logic valid;
    logic [31:0] addr;
    logic [31:0] data_mem;
    logic [6:0] pd_reg;
    logic [4:0] rob_reg;
    logic load_en;
    
    // LSQ
    logic store_wb;
    lsq lsq_out;
    logic lsq_full;
    
    always_comb begin
        // L-type and S-type instructions
        if (data_in.Opcode == 7'b0000011) begin
            addr = ps1_data + data_in.imm;
        end else begin
            addr = '0;
        end
    end    
    
    always_ff @(posedge clk or posedge reset) begin
        if (reset) begin
            load_en <= 1'b0;
            pd_reg     <= '0;
            rob_reg    <= '0;
        end else begin
            if (mispredict) begin
                load_en <= 1'b0;
            end else begin
                if (issued && data_in.Opcode == 7'b0000011 && !load_en) begin
                    load_en <= 1'b1;
                    pd_reg     <= data_in.pd;
                    rob_reg    <= data_in.rob_index;
                end

                // Clear when memory returns valid data
                if (valid && load_en) begin
                    load_en <= 1'b0;
                end
            end
        end
    end
    
    always_comb begin   
        data_out.fu_mem_ready = 1'b1;
        data_out.fu_mem_done  = 1'b0;
        data_out.p_mem = '0;
        data_out.rob_fu_mem = '0;
        data_out.data = '0;
        
        
        if (load_en) begin
            data_out.fu_mem_ready = 1'b0;
        end 
        
        // stall if we're full when store
        if (data_in.Opcode == 7'b0100011 && lsq_full) begin
            data_out.fu_mem_ready = 1'b0;
        end
        
        if (mispredict) begin
            automatic logic [4:0] ptr = (mispredict_tag == 15) ? 0 : mispredict_tag + 1;
            for (logic [4:0] i = ptr; i != curr_rob_tag; i=(i==15)?0:i+1) begin
                if (i == data_in.rob_index) begin
                    data_out.p_mem = '0;
                    data_out.rob_fu_mem = '0;
                    data_out.data = '0;
                    data_out.fu_mem_ready = 1'b1;
                    data_out.fu_mem_done = 1'b0;
                end
            end
        end else begin
            if (issued) begin
                if (data_in.Opcode == 7'b0100011 && !lsq_full) begin // sw
                    data_out.fu_mem_ready = 1'b1;
                    data_out.fu_mem_done = 1'b1;
                    data_out.rob_fu_mem = data_in.rob_index;
                end else if (data_in.Opcode == 7'b0000011 && !load_en) begin // lw
                    data_out.fu_mem_ready = 1'b0;
                    data_out.fu_mem_done = 1'b0;
                    data_out.p_mem = data_in.pd;
                    data_out.rob_fu_mem = data_in.rob_index;
                end
            end
            if (valid && load_en) begin
                data_out.fu_mem_ready = 1'b1;      // free again
                data_out.fu_mem_done  = 1'b1;
                data_out.p_mem        = pd_reg;
                data_out.rob_fu_mem   = rob_reg;
                data_out.data         = data_mem;
            end
        end
    end
    
    lsq u_lsq (
        .clk(clk),
        .reset(reset),
        
        .ps1_data(ps1_data),
        .imm_in(data_in.imm),
        
        // From PRF
        .ps2_data(ps2_data),
        
        .issued(issued),
        .data_in(data_in),
        
        // From ROB
        .retired(retired),
        .rob_head(rob_head),
        .store_wb(store_wb),
        .data_out(lsq_out),
        .full(lsq_full) 
    );
    
    data_memory u_dmem (
        .clk(clk),
        .reset(reset),
        
        .addr(addr),
        .issued(issued),
        .Opcode(data_in.Opcode),
        .func3(data_in.func3),
        
        // From LSQ for S-type
        .store_wb(store_wb),
        .lsq_in(lsq_out),
        
        .data_out(data_mem),
        .valid(valid)
    );
    
endmodule
